
module Quasi6502
   (input  wire         reset,
    output wire         ready,
    input  wire         clk,
    input  wire         irq,
    input  wire         nmi,
    output wire         sync,
    output wire         busRequestWrite,
    output wire [15:0]  busRqAddress,
    input  wire  [7:0]  busDataIn,
    output wire  [7:0]  busDataOut);

    // STUB.
endmodule

